'`timescale 1ns/1ns
'`include "first.v"

module fir (
    ports
);
    
endmodule